.title 4th Order Butterworth LPF
.include "~/Documents/SPICE/TL074.lib"
.save all

XU1 /b /c +3.3V -3V3 /c TL074
C4 v_out /d 680p
R4 /d /e 1k
R3 /c /d 1.3k
C3 0 /e 100p
XU3 /e v_out +3.3V -3V3 v_out TL074
R2 /a /b 2.2k
R1 v_in /a 3k
V1 -3V3 0 DC -3.3 
C1 0 /b 100p
V3 +3.3V 0 DC 3.3 
V2 v_in 0 DC 500m SIN( 500m 500m 1k 0 0 0 500m ) AC 500m 
C2 /c /a 120p

.control
ac dec 100k 10 100Meg
* settype decibel out
* plot vdb(v_out) xlimit 1 100Meg ylabel 'Magnitude (dB)'
* settype phase out
* plot cph(v_out) xlimit 1 100Meg ylabel 'phase (rad/s)'
* let outd = 180/PI*cph(v_out)
* settype phase outd
* plot outd xlimit 1 100Meg ylabel 'phase (degrees)'
wrdata vdb_data vdb(v_out)
wrdata vp_data vp(v_out)
quit
.endc

.end

